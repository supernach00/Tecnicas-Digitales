LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ConvGRAYaBIN IS 
	PORT(
		
		GRAY_IN : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		BIN_OUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	
	);
	
END ConvGRAYaBIN;

ARCHITECTURE ARCH1 OF ConvGRAYaBIN IS


	TYPE FORMATO_ROM IS ARRAY (0 TO 7) OF STD_LOGIC_VECTOR(2 DOWNTO 0);
	CONSTANT ROM : FORMATO_ROM := (
	
	"000",   -- GRAY 000
	"001",   -- GRAY 001
	"011",   -- GRAY 010
	"010",   -- GRAY 011
	"111",   -- GRAY 100
	"110",   -- GRAY 101
	"100",   -- GRAY 110
	"101"   -- GRAY 111
	
	);
	

BEGIN

	BIN_OUT <= ROM(TO_INTEGER(UNSIGNED(GRAY_IN)));
	
END ARCHITECTURE;