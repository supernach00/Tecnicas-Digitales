library verilog;
use verilog.vl_types.all;
entity flipflops_vlg_vec_tst is
end flipflops_vlg_vec_tst;
