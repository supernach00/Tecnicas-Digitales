library verilog;
use verilog.vl_types.all;
entity nacho_vlg_vec_tst is
end nacho_vlg_vec_tst;
