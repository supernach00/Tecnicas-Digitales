library verilog;
use verilog.vl_types.all;
entity proceso2_vlg_vec_tst is
end proceso2_vlg_vec_tst;
